library verilog;
use verilog.vl_types.all;
entity test_vlg_tst is
end test_vlg_tst;
